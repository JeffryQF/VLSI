*** SPICE deck for cell Or-Or-And-Inv{sch} from library Tarea_2_VLSI
*** Created on lun oct 05, 2015 14:06:41
*** Last revised on lun oct 12, 2015 18:07:36
*** Written on lun oct 12, 2015 19:06:28 by Electric VLSI Design System, version 9.06
*** Layout tech: mocmos, foundry MOSIS
*** UC SPICE *** , MIN_RESIST 4.0, MIN_CAPAC 0.1FF

.global gnd vdd

*** TOP LEVEL CELL: Or-Or-And-Inv{sch}
Mnmos@0 _F A net@13 gnd NMOS L=0.6U W=6.666U
Mnmos@1 _F B net@13 gnd NMOS L=0.6U W=6.666U
Mnmos@2 net@13 C gnd gnd NMOS L=0.6U W=6.666U
Mnmos@3 net@13 D gnd gnd NMOS L=0.6U W=6.666U
Mpmos@0 vdd A net@3 vdd PMOS L=0.6U W=11.328U
Mpmos@1 vdd D net@67 vdd PMOS L=0.6U W=11.328U
Mpmos@2 net@3 B _F vdd PMOS L=0.6U W=11.328U
Mpmos@3 net@67 C _F vdd PMOS L=0.6U W=11.328U

* Spice Code nodes in cell cell 'Or-Or-And-Inv{sch}'
Vdd vdd 0 DC 3.3
Vin A 0 PULSE(0 3.3 0 0 0 1n 2n 2)
.tran 1n 4n
.include C:\Users\Francis\Desktop\Electric (VLSI)\Mosis_5.txt
.END
