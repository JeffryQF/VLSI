*** SPICE deck for cell Inversor_dinamico{sch} from library Tarea_1_VLSI
*** Created on mar sep 01, 2015 23:17:26
*** Last revised on sáb sep 12, 2015 09:45:48
*** Written on sáb sep 12, 2015 09:45:56 by Electric VLSI Design System, version 9.06
*** Layout tech: mocmos, foundry MOSIS
*** UC SPICE *** , MIN_RESIST 4.0, MIN_CAPAC 0.1FF

.global gnd vdd

*** TOP LEVEL CELL: Inversor_dinamico{sch}
Mnmos@0 out in gnd gnd N L=0.18U W=1.08U
Mpmos@0 vdd in out vdd P L=0.18U W=2.16U

* Spice Code nodes in cell cell 'Inversor_dinamico{sch}'
vdd vdd 0 DC 3.3
Vin in 0 DC 0
.dc Vin 0 3.3 1m
.include C:\Users\Francis\Desktop\Electric (VLSI)\C5_models.txt
.END
